

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity noisy_signal is
    Port ( 
        addr : in unsigned(9 downto 0);
        data_out : out signed(15 downto 0)
    );
end noisy_signal;

architecture Behaviroal of noisy_signal is 

    
type signal_value is array (0 to 999) of signed(15 downto 0);

-- Declare the constant using the defined type
constant signal_array : signal_value := (
    "0001000010101101",
    "0000101011101101",
    "1111101110010111",
    "0001101011100100",
    "0010111001010011",
    "0011001011110011",
    "0011111101001100",
    "0011010001010011",
    "0011001110110100",
    "0100010101001001",
    "0100100100110110",
    "0100110010111111",
    "0100000111000111",
    "0101100010010000",
    "0110001010100010",
    "0011010110101010",
    "0100110011001001",
    "0100000000111101",
    "0100001110010111",
    "0100000100000101",
    "0100101110111110",
    "0100000001010001",
    "0011100111011101",
    "0011111111100000",
    "0011111011100001",
    "0011111010000110",
    "0011100000100110",
    "0011111000100011",
    "0011110111100110",
    "0011110100000110",
    "0101101001011100",
    "0101010001011110",
    "0100101111000100",
    "0101011100110101",
    "0100100001111110",
    "0101000111010001",
    "0100100110001011",
    "0100010001011000",
    "0100000101011100",
    "0110010001001011",
    "0100111100001100",
    "0100111110111111",
    "0100011110100010",
    "0100111001001001",
    "0101110000111101",
    "0100011000110101",
    "0011100111110001",
    "0011000000111100",
    "0010100101011001",
    "0001101110011000",
    "0010011100101100",
    "0010100101001101",
    "0001110110011100",
    "0001010001000001",
    "0001110100000001",
    "0000101000000100",
    "0001001011001100",
    "1111101100100010",
    "0000011110100000",
    "1111110010001010",
    "0000011101110010",
    "0000001111110111",
    "0000101001000100",
    "0000010111010011",
    "1111110011000111",
    "0000011111110000",
    "0001000001010011",
    "0001011110011001",
    "0000101110001011",
    "0001001001101000",
    "0001011110110011",
    "0001111001101000",
    "0010010000111000",
    "0011000011111110",
    "0001101011101100",
    "0011100111110000",
    "0010000010001010",
    "0010101110000110",
    "0001100111110110",
    "0010100001100010",
    "0011001100101010",
    "0010101110110011",
    "0010000101111000",
    "0001111000000001",
    "0001000110001000",
    "0001011000101101",
    "0001110000110111",
    "0000110110100010",
    "0001001100100001",
    "0001101010100101",
    "0001010001110011",
    "0001010100111101",
    "0000100111010111",
    "0001011010111111",
    "0001010111010100",
    "0010010000001011",
    "0000100010011001",
    "0000111011011111",
    "0001001111101001",
    "0001101011000010",
    "0001011001110110",
    "0011011011111110",
    "0011000111001011",
    "0010111011000000",
    "0010100010111111",
    "0011001000111001",
    "0010011111110011",
    "0001101010110001",
    "0011010101010100",
    "0011101101110100",
    "0010010110101101",
    "0010100010001010",
    "0001010001111101",
    "0001100101111011",
    "0001010000111111",
    "0000011000111100",
    "1111011110111010",
    "1111111111010010",
    "0000000010101011",
    "1110110111100011",
    "1101011101011000",
    "1101101101010011",
    "1100101110111000",
    "1100101100000110",
    "1011110101000111",
    "1100111110011100",
    "1011010010010101",
    "1010001110000111",
    "1010111101111111",
    "1100111010001111",
    "1011111110110110",
    "1010110111110001",
    "1011011110010011",
    "1011101000000010",
    "1010100101001000",
    "1011101011010001",
    "1011001101011011",
    "1011110110011011",
    "1011111100101110",
    "1001110010110010",
    "1011000111110100",
    "1011011001100010",
    "1100010010101101",
    "1010001101110001",
    "1011010101001110",
    "1010000111100010",
    "1011000100011001",
    "1011010011111011",
    "1010100101100100",
    "1010000111000100",
    "1001111101110011",
    "1000101101111111",
    "1010001100111010",
    "1000011001010110",
    "1000111111100101",
    "1001100101100000",
    "1000000101110011",
    "1000011110101110",
    "1001100101111001",
    "1001111011111100",
    "1010011110011100",
    "1010111110100110",
    "1011001001100001",
    "1011001000010000",
    "1011000011100110",
    "1011110010100110",
    "1100101111001101",
    "1101010001100010",
    "1101000011110110",
    "1101110100100001",
    "1110110001111100",
    "1111000001111100",
    "1111011110110010",
    "1111010010000010",
    "1111110010100110",
    "1111101011110010",
    "1111010000100000",
    "0000111010101011",
    "0000011011111110",
    "0000000011000110",
    "1111101110101000",
    "0000101101010111",
    "0001100110100001",
    "1111100001111110",
    "0000111101111001",
    "0001001001011000",
    "1111011100000101",
    "0000001000111101",
    "1111110111000111",
    "0001000000011011",
    "0000000110100101",
    "0000100001111100",
    "0000010110011010",
    "0000100001011100",
    "1111101010011000",
    "1111111011011001",
    "0000011010011110",
    "0000101100011100",
    "0000110001110000",
    "0001011001001011",
    "0001111110010101",
    "0000100110011111",
    "0000111001110001",
    "0010100011100001",
    "0010100011111111",
    "0011000000111010",
    "0001011010010011",
    "0010101001000000",
    "0010110111101110",
    "0001101100010000",
    "0010000100110000",
    "0011001000000000",
    "0001110011111110",
    "0001100010010110",
    "0001010111011111",
    "0000110110001010",
    "0000100010000011",
    "0000000001110101",
    "0000100000000111",
    "0000011111110001",
    "1110110010011100",
    "0000010000010100",
    "0000000011101100",
    "1110001100101110",
    "1111000101100010",
    "1111100110010010",
    "0000001110010101",
    "1110110010111100",
    "1111011011100111",
    "0000110011001010",
    "0000000110000001",
    "1111110000000111",
    "0001010000111111",
    "0001010000010110",
    "0001110110001000",
    "0001111110000100",
    "0010010101101000",
    "0010011011010110",
    "0011000110101001",
    "0011111011110101",
    "0011011111110011",
    "0010000010000111",
    "0010111001010111",
    "0101001000011110",
    "0100000001110100",
    "0100010001111011",
    "0010111110101100",
    "0011000101001000",
    "0100010110010111",
    "0100000110001000",
    "0100001011011010",
    "0100010101010111",
    "0100000100101001",
    "0010111011111001",
    "0100100011010000",
    "0011000101110100",
    "0100000011101100",
    "0010110111100011",
    "0010111111011110",
    "0011111101000000",
    "0100000010000100",
    "0011100110010111",
    "0101101100101100",
    "0100010101101010",
    "0101110001000001",
    "0110111011000000",
    "0110010000000000",
    "0101100011000111",
    "0111000001001100",
    "0110110011001010",
    "0110111100101011",
    "0110111001010101",
    "0110000010001100",
    "0111001110010110",
    "0101011011111101",
    "0110111011000001",
    "0101101010000110",
    "0110001100011000",
    "0110001010001101",
    "0101000000010000",
    "0110101010010011",
    "0100000011101110",
    "0100010000100011",
    "0011011000111001",
    "0011110010110011",
    "0000111111011001",
    "0010000100110010",
    "0000111111101011",
    "0010010111011001",
    "1111100110101101",
    "0000010100101010",
    "0001110110111111",
    "1111001101110011",
    "1111101101001110",
    "1111110010100101",
    "1110101101100001",
    "1110111011100010",
    "1110101100001001",
    "1110111101110110",
    "1110010000010000",
    "1110110101100011",
    "1101111000000111",
    "1110100011101001",
    "1101010011000001",
    "1101011010101000",
    "1110111101000000",
    "1110111001000101",
    "1110101101101000",
    "1101111111001001",
    "1101001111110011",
    "1101100000001000",
    "1100111100111010",
    "1110100011100100",
    "1100011001111111",
    "1101100100111100",
    "1010111100111100",
    "1100011000011010",
    "1011100111000111",
    "1011101011011000",
    "1010100011011101",
    "1010011111101101",
    "1010100111110000",
    "1011111010110100",
    "1010110001000010",
    "1001010000100010",
    "1010100110000000",
    "1010111000100110",
    "1010111000101100",
    "1011011010110111",
    "1011101110110110",
    "1011011010111111",
    "1100100010001100",
    "1100000011000011",
    "1011011000000001",
    "1100110000000000",
    "1100111000001101",
    "1101011001101111",
    "1110011001000101",
    "1110101100011011",
    "1110111001101011",
    "1110100100000010",
    "1110111111000110",
    "0000101101110000",
    "1111110010110010",
    "1110111010111101",
    "0000001100110101",
    "1110011110001011",
    "1110000011100110",
    "1110111010010000",
    "1110100110011001",
    "1110110100000110",
    "1110110100001011",
    "1101000100000100",
    "1110010000101000",
    "1101101000000111",
    "1101010001101110",
    "1100011011001111",
    "1101011010101010",
    "1101010101110000",
    "1101010001111110",
    "1100001110001101",
    "1101110010000101",
    "1111000110001011",
    "1100100100110010",
    "1110000111100010",
    "1101010000011000",
    "1110001001000011",
    "1110001011100010",
    "1110110000100111",
    "1110111101011110",
    "1111100000110100",
    "1110011110110001",
    "1111011100100001",
    "1110111100100100",
    "1111000000111100",
    "1111110100000101",
    "1110110100001010",
    "1110001110011110",
    "1110100001110011",
    "1101011001101011",
    "1101111010011100",
    "1100000001000100",
    "1100110101011011",
    "1011100100100000",
    "1011101011011000",
    "1101000101000000",
    "1010111011100101",
    "1010111010000110",
    "1011010110111001",
    "1100010110000101",
    "1010000011110011",
    "1011001101101100",
    "1011111011001000",
    "1011001100111111",
    "1011000101010001",
    "1010101100001111",
    "1011110110011100",
    "1011010010001110",
    "1101101111011001",
    "1101010010000101",
    "1100001001110001",
    "1101011101011100",
    "1110111001011111",
    "1111101000000110",
    "0000001000000001",
    "1111111100111111",
    "0001000010111000",
    "1111100110011100",
    "0001010101000010",
    "0001111011110011",
    "0000111000011100",
    "0000110100011010",
    "0010111011001001",
    "0001011011100101",
    "0001010101110000",
    "0010001110011000",
    "0001111011111000",
    "0000111110101101",
    "0010101000110100",
    "0010001010101001",
    "0001110000010111",
    "0010001100000000",
    "0010110001010000",
    "0001100011010110",
    "0001010101000011",
    "0010010100111100",
    "0011001101110101",
    "0011000100010001",
    "0100111101101111",
    "0100010011010111",
    "0101001011011001",
    "0011011100110110",
    "0101001111111101",
    "0101100011000100",
    "0101010100001010",
    "0110010010000001",
    "0110011101000010",
    "0110100101110010",
    "0110011101010100",
    "0111001001100000",
    "0111100000010110",
    "0111111111111111",
    "0110101101000010",
    "0111011000110100",
    "0110100110001001",
    "0111011010101111",
    "0110110111101001",
    "0101011101001111",
    "0101111010010001",
    "0101110011011100",
    "0101010101000100",
    "0100111000001101",
    "0011111011111001",
    "0101001000111110",
    "0011101010100010",
    "0011011111100110",
    "0011101100101010",
    "0011101111010110",
    "0001110011100110",
    "0010011010011101",
    "0010101010000111",
    "0001100000111001",
    "0001110110110100",
    "0001110001001000",
    "0000110111010001",
    "0000110011100101",
    "0011001001000111",
    "0001011110011110",
    "0001010101100011",
    "0010000111100001",
    "0010010100001001",
    "0010001010000011",
    "0010100011100011",
    "0001111111000110",
    "0010001110011000",
    "0010000000010111",
    "0000101111011101",
    "1111010000000011",
    "0001100011111100",
    "0001000010101011",
    "0001000101111000",
    "0000000110111010",
    "1111011011111100",
    "1111110100010100",
    "1111000100100010",
    "1110011001000101",
    "1110001010101001",
    "1101110010111101",
    "1110110001000010",
    "1110010100000101",
    "1110010001010000",
    "1110100100000100",
    "1101101101000001",
    "1110110111110110",
    "1110001101011101",
    "1110101010101000",
    "1111001010001010",
    "1110100110000110",
    "1111000111010110",
    "0000101100001101",
    "0000001010010111",
    "0000000010000010",
    "0000101010100000",
    "0001000000100110",
    "0000110111110101",
    "0000001011001101",
    "0001100100111000",
    "0000101101111111",
    "0000110000011001",
    "0001010101000101",
    "0010110111010011",
    "0010000111100011",
    "0010000010101100",
    "0000110010001110",
    "0001011110110001",
    "0001010100111010",
    "0000110110001000",
    "0000010100000000",
    "1111011100110000",
    "0000110100001010",
    "1110000011010100",
    "1110101110100011",
    "1111000001101100",
    "1110111111010111",
    "1110001111001110",
    "1110110111001010",
    "1110110010101111",
    "1110001000011011",
    "1110100101111100",
    "1101100100000000",
    "1110110101000111",
    "1110101001111111",
    "1110111111000111",
    "1110001111001011",
    "1100111101100011",
    "1110000101111011",
    "1101101111010001",
    "1110101001010000",
    "1101111101110111",
    "1110001011010001",
    "1110011100011100",
    "1110100001101010",
    "1110010010101100",
    "1101010011110000",
    "1100111101100110",
    "1100001100101000",
    "1101100111010011",
    "1100001011010011",
    "1100100011100111",
    "1100010111011010",
    "1011010110010111",
    "1011011111110010",
    "1010000110010000",
    "1000001110110111",
    "1001000010001111",
    "1000110010011110",
    "1000001011101111",
    "1000010100101011",
    "1010000111100000",
    "1000010001010100",
    "1001010011101110",
    "1001001100101110",
    "1000010100100100",
    "1000110100110001",
    "1000010111101011",
    "1000111100100111",
    "1010001100111111",
    "1001111010000000",
    "1011010000010000",
    "1010111011111001",
    "1010111011001011",
    "1100010100110000",
    "1100010100101011",
    "1100011110000111",
    "1100001111110000",
    "1100111000111011",
    "1110010100101010",
    "1101001011101010",
    "1101000000001000",
    "1110011101101100",
    "1101110000010110",
    "1110000010011010",
    "1110110101101011",
    "1101100100011011",
    "1110110110001111",
    "1110011001010000",
    "1111001010101101",
    "1101101011100111",
    "1101010110110100",
    "1110100000001010",
    "1111101101111010",
    "1110111111101100",
    "1111000110100010",
    "1111000101010111",
    "0000100101101110",
    "0000111010111011",
    "0000110000110111",
    "0001110101111011",
    "0011001000001001",
    "0010010011001101",
    "0010000010011110",
    "0011010010100011",
    "0011110101111110",
    "0100000010011101",
    "0100000010001011",
    "0100000100010011",
    "0011110000010101",
    "0101000101101111",
    "0100110011111100",
    "0101000111001110",
    "0100110001011111",
    "0100101011001111",
    "0011111100110011",
    "0100000011000101",
    "0100001011111111",
    "0011111011101001",
    "0100000001111101",
    "0011010111110011",
    "0010001101011101",
    "0001111101111111",
    "0011000010111100",
    "0001100010101000",
    "0001101000111011",
    "0001100001111111",
    "0001100100111000",
    "0001001010100001",
    "0001100001000110",
    "0000001110100010",
    "0001111011100100",
    "0000011100010001",
    "0010000011001110",
    "0001110111001100",
    "0001100111000011",
    "0001101111001011",
    "0010000100100110",
    "0001110110000101",
    "0010011011100110",
    "0010010000001111",
    "0010101000000010",
    "0011111010001000",
    "0001011110100110",
    "0001110111110000",
    "0010011111000011",
    "0010001100100001",
    "0011011000001011",
    "0010001001100000",
    "0001111111011101",
    "0010100011111111",
    "0001100100010100",
    "0001011011110001",
    "0001011100000000",
    "0000111111110111",
    "0001001000001010",
    "0000000101000011",
    "0001001010101100",
    "0000010110100010",
    "0000100100111010",
    "0000111101110011",
    "0001100011111100",
    "0001010010111001",
    "0000110010101100",
    "0001011011100011",
    "0001101100000100",
    "0001101111011100",
    "0011010010001100",
    "0011000110010011",
    "0011100111100010",
    "0100000010100101",
    "0011011000000001",
    "0011111011111011",
    "0100100010101101",
    "0101011100110101",
    "0100101010110100",
    "0110000101010001",
    "0101101101110101",
    "0110000101001111",
    "0101000100001001",
    "0110110100111010",
    "0101101110011100",
    "0100111010111111",
    "0110000110110000",
    "0100110001101000",
    "0100001001010000",
    "0101100011010001",
    "0011101101000110",
    "0011100111010011",
    "0100000101011010",
    "0010101110110110",
    "0011000011001010",
    "0011111010000010",
    "0000110111110010",
    "0011000010111101",
    "0001101011011110",
    "0001111000000110",
    "0001101011010110",
    "0010000101111101",
    "0001011111111101",
    "0001110001001101",
    "0000101111101111",
    "0001010001101111",
    "0001001110101010",
    "0001001010011110",
    "0001011111010101",
    "0010000011000101",
    "0001000110110110",
    "0010011101000100",
    "0000010000001011",
    "0001001011001011",
    "1111111011000000",
    "0000110010000001",
    "1111111100011001",
    "1110101110000100",
    "1110101110110000",
    "1110011011010110",
    "1110100011100001",
    "1101011101111000",
    "1101100110110111",
    "1100110011011111",
    "1011010110011101",
    "1010111101111001",
    "1011110100001100",
    "1010010001110011",
    "1011001101011000",
    "1011001111001000",
    "1001011110101110",
    "1001111110111001",
    "1010010010100100",
    "1001110000000011",
    "1001110011011100",
    "1001011001011110",
    "1001001100000011",
    "1010010100100101",
    "1001010110101101",
    "1001011111011101",
    "1010001011010111",
    "1011100000000010",
    "1011001101110010",
    "1100000001001110",
    "1011111011110101",
    "1011110111100110",
    "1100000100011011",
    "1100110001110100",
    "1011000111000101",
    "1100101011101011",
    "1100011000001110",
    "1011101100001101",
    "1100001010100000",
    "1100111011101100",
    "1100100100100000",
    "1011010100010010",
    "1100100100100001",
    "1100100000001011",
    "1011011111111000",
    "1101010010011011",
    "1011111100110010",
    "1011001010110110",
    "1010110101001100",
    "1100010100010110",
    "1100101111101001",
    "1100000011000111",
    "1101000000011101",
    "1101110111101001",
    "1110110010110100",
    "1101110001001011",
    "1101010010000010",
    "1110001111000001",
    "1110000001001101",
    "1111110001001111",
    "1111110111000100",
    "1111110010011000",
    "1111001101010000",
    "0000001010100001",
    "0000110101111111",
    "0000011000011001",
    "0001011010010110",
    "0001111111111111",
    "0000101000000100",
    "0000010010000001",
    "0001001111101100",
    "0000010000101100",
    "0001011111100100",
    "0000001000001010",
    "1111110001111001",
    "1110101010101111",
    "1111110000011100",
    "1111011110011000",
    "1110011010001111",
    "1110011110010110",
    "1110110001100001",
    "1101111011100001",
    "1110101101000010",
    "1110000111100000",
    "1101010001000000",
    "1110000110000101",
    "1101000001000011",
    "1100100111000101",
    "1110010111110000",
    "1110001111000100",
    "1110011110110010",
    "1101000110010010",
    "1101010110111010",
    "1111000110111111",
    "1111000000001100",
    "1110011110111000",
    "1110000011001001",
    "1110010001100101",
    "0000110101011100",
    "1110101000111111",
    "0000101111011110",
    "1111000001011110",
    "1111100010000001",
    "1111000010100111",
    "0000001100100111",
    "1110111101100110",
    "1111010001101000",
    "1110111010110001",
    "1111011111110111",
    "1111011101011010",
    "0000000000101001",
    "1111110010101101",
    "1110101101100000",
    "1110111110001001",
    "1110101000000011",
    "1111100110001011",
    "0000010101000001",
    "1111111110110100",
    "0000011011001001",
    "1111110001110111",
    "0001000110000011",
    "0001011001001001",
    "0001100001100101",
    "0010000111000011",
    "0010111100110101",
    "0010001001000011",
    "0011100000010100",
    "0011110111101110",
    "0011100101010001",
    "0100111010110011",
    "0101011100101101",
    "0100100000000111",
    "0110010111000100",
    "0101010000100101",
    "0110100011100111",
    "0110000011101010",
    "0110010111111110",
    "0111101000101000",
    "0110100100000100",
    "0110110011011001",
    "0110011010111100",
    "0110000111101100",
    "0110011111001001",
    "0110000011110111",
    "0101010010100100",
    "0110010101100001",
    "0101000010001001",
    "0100011111001100",
    "0100111010110000",
    "0110000101001010",
    "0100011111111101",
    "0100101011100010",
    "0101010011000001",
    "0100101010110011",
    "0101110011110011",
    "0100101010101111",
    "0100000111100011",
    "0011110001100011",
    "0100010100010000",
    "0100101111001110",
    "0100000000110101",
    "0101000110000100",
    "0100101001111101",
    "0100110111100000",
    "0100011100111111",
    "0011111100110100",
    "0011110111011000",
    "0100000110011001",
    "0011001010100101",
    "0010001010110111",
    "0001110010101101",
    "0010000110101110",
    "0010000100111001",
    "0001010101010011",
    "0001101101000010",
    "1111111101011100",
    "0000100000100111",
    "1110111100001011",
    "1111011001101101",
    "1111001100111100",
    "1110110011001111",
    "1101011001110101",
    "1110000010001111",
    "1110001011111001",
    "1101010101010110",
    "1101101000001011",
    "1101110111011001",
    "1101000011011000",
    "1011100110011001",
    "1100111001011100",
    "1011111100111101",
    "1110000110100000",
    "1101100111010111",
    "1100110000101101",
    "1101001001101101",
    "1110000001001111",
    "1110111010100010",
    "1110000001111010",
    "1110010101000010",
    "1111001101100001",
    "1111000100010001",
    "1110010110101011",
    "1110111101010100",
    "1111011011111011",
    "1110011110001001",
    "1110111101001010",
    "1110100111110100",
    "1101111101010010",
    "1101111110110000",
    "1110110100101010",
    "1110000011010111",
    "1110000001010010",
    "1101111110010011",
    "1101101001111110",
    "1101111010001001",
    "1101010001110001",
    "1101100110110010",
    "1101110100000100",
    "1101110110111011",
    "1110010111010110",
    "1101111101100101",
    "1110011100100000",
    "1110101000010001",
    "1101110001011101",
    "1110010011011000",
    "1111010001010011",
    "0000110111011010",
    "1110101011011101",
    "1111111001101110",
    "1111010111110111",
    "1111011011000100",
    "0000010010011010",
    "1111100011111011",
    "0001000101011011",
    "1111001101101101",
    "1111111010101000",
    "0000010010001101",
    "1111001001000100",
    "1111000011101010",
    "1110100111110010",
    "1101111001000110",
    "1110101100111010",
    "1101100100000001",
    "1110101000101100",
    "1100110100110110",
    "1011111110101111",
    "1011111101000111",
    "1011001101101000",
    "1100001011101110",
    "1010110110100010",
    "1010100010111111",
    "1010001100101100",
    "1011001110110000",
    "1010101010000011",
    "1011000010010000",
    "1010101000000100",
    "1100001001010111",
    "1010001111011000",
    "1011001110101001",
    "1010101010110010",
    "1010110001100010",
    "1011011101011010",
    "1011010111100110",
    "1100001101100111",
    "1011110100111110",
    "1011101110110011",
    "1100101101101000",
    "1100000110110110",
    "1011110000101011",
    "1100000110100010",
    "1100010101001100",
    "1011001100000010",
    "1100100001011001",
    "1011111111001110",
    "1010110000000101",
    "1011001111111001",
    "1100011010001010",
    "1011101101011111",
    "1100101001101101",
    "1011000111111011",
    "1100000111000010",
    "1100000100100001",
    "1011011011010101",
    "1011110101100011",
    "1101000111111111",
    "1101000111001011",
    "1100101100100000",
    "1101100101110100",
    "1110011011100000",
    "1110001000010110",
    "1110010111010000",
    "1111110011001010"

);

begin
    
    data_out <= signal_array(to_integer(addr));


end Behaviroal;