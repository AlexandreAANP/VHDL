library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity filter_rom is
    Port ( 
        addr : in std_logic_vector(5 downto 0);
        data_out : out std_logic_vector(15 downto 0)
    );
end filter_rom;

architecture Behaviroal of filter_rom is 

    
type coeff_array is array (0 to 50) of signed(15 downto 0);

-- Declare the constant using the defined type
constant coeffs : coeff_array := (
    "0000000000000000",
    "0000000000000001",
    "0000000000000010",
    "0000000000000011",
    "0000000000000100",
    "0000000000000101",
    "0000000000000110",
    "0000000000000111",
    "0000000000001000",
    "0000000000001001",
    "0000000000001010",
    "0000000000001011",
    "0000000000001100",
    "0000000000001101",
    "0000000000001110",
    "0000000000001111",
    "0000000000010000",
    "0000000000010001",
    "0000000000010010",
    "0000000000010011",
    "0000000000010100",
    "0000000000010101",
    "0000000000010110",
    "0000000000010111",
    "0000000000011000",
    "0000000000011001",
    "0000000000011010",
    "0000000000011011",
    "0000000000011100",
    "0000000000011101",
    "0000000000011110",
    "0000000000011111",
    "0000000000100000",
    "0000000000100001",
    "0000000000100010",
    "0000000000100011",
    "0000000000100100",
    "0000000000100101",
    "0000000000100110",
    "0000000000100111",
    "0000000000101000",
    "0000000000101001",
    "0000000000101010",
    "0000000000101011",
    "0000000000101100",
    "0000000000101101",
    "0000000000101110",
    "0000000000101111",
    "0000000000110000",
    "0000000000110001",
    "0000000000110001"
);

begin
    
    data_out <= std_logic_vector(coeffs(to_integer(unsigned(addr))));


end Behaviroal;